// module imem (
// 	a,
// 	instr_addr
// );
// 	// memory position to access/index
// 	input wire [31:0] a;
// 	// read data reg
// 	output wire [31:0] instr_addr;
	
// 	// access RAM 'a' position
// 	// assign instr_addr = a[31:2];

// endmodule

module imem (
	a,
	rd
);
	// memory position to access/index
	input wire [31:0] a;
	// read data reg
	output wire [31:0] rd;
	
	wire [31:0] RAM [3:0];

	assign RAM[0] = 32'h00500113;
	assign RAM[1] = 32'h00c00193;
	assign RAM[2] = 32'h01e00113;
	assign RAM[3] = 32'h02202423;
		
	// access RAM 'a' position
	assign rd = RAM[a[31:2]];

endmodule


//{
//32'h00500113,
//32'h00c00193
//};
// 32'hff718393,
// 32'h0023e233,
// 32'h0041f2b3,
// 32'h004282b3,
// 32'h02728863,
// 32'h0041a233,
// 32'h00020463,
// 32'h00000293,
// 32'h0023a233,
// 32'h005203b3,
// 32'h402383b3,
// 32'h0471aa23,
// 32'h06002103,
// 32'h005104b3,
// 32'h008001ef,
// 32'h00100113,
// 32'h00910133,
// 32'h0221a023,
// 32'h000010b7,
// 32'h06102423,
// 32'h00001097,
// 32'h06102623,
// 32'h06100193,
// 32'h00f180e7,
// 32'h00100193,
// 32'h00200193,
// 32'h06102823,
// 32'hfff00113,
// 32'h00200193,
// 32'h00312233,
// 32'h06402a23,
// 32'hfff00113,
// 32'h00200193,
// 32'h00313233,
// 32'h06402c23,
// 32'h00900093,
// 32'h00900113,
// 32'h00208463,
// 32'h00800093,
// 32'h06102e23,
// 32'h00900093,
// 32'h00a00113,
// 32'h00209463,
// 32'h00800093,
// 32'h08102023,
// 32'hfff00093,
// 32'h00100113,
// 32'h0020c463,
// 32'h00800093,
// 32'h08102223,
// 32'h00100093,
// 32'hfff00113,
// 32'h0020d463,
// 32'h00800093,
// 32'h08102423,
// 32'h00100093,
// 32'hfff00113,
// 32'h0020e463,
// 32'h00800093,
// 32'h08102623,
// 32'hfff00093,
// 32'h00100113,
// 32'h0020f463,
// 32'h00800093,
// 32'h08102823,
// 32'h05400093,
// 32'h0aa00113,
// 32'h0020c1b3,
// 32'h08302a23,
// 32'h09800093,
// 32'h0260c193,
// 32'h08302c23,
// 32'h0720e193,
// 32'h08302e23,
// 32'h06a0f193,
// 32'h0a302023,
// 32'hfff0a193,
// 32'h0a302223,
// 32'hfff0b193,
// 32'h0a302623,
// 32'hfb300093,
// 32'h00109193,
// 32'h06302223,
// 32'h0010d193,
// 32'h06302423,
// 32'h4010d193,
// 32'h06302623,
// 32'h00100113,
// 32'h002091b3,
// 32'h06302823,
// 32'h0020d1b3,
// 32'h06302a23,
// 32'h4020d1b3,
// 32'h06302c23,
// 32'haa0bc0b7,
// 32'h0dd08093,
// 32'h06102023,
// 32'h06000103,
// 32'h0a202023,
// 32'h06100103,
// 32'h0a202223,
// 32'h06200103,
// 32'h0a202423,
// 32'h06300103,
// 32'h0a202623,
// 32'h06001103,
// 32'h0a202823,
// 32'h06101103,
// 32'h0a202a23,
// 32'h06201103,
// 32'h0a202c23,
// 32'h06301103,
// 32'h0a202e23,
// 32'h06004103,
// 32'h06202223,
// 32'h06104103,
// 32'h06202423,
// 32'h06204103,
// 32'h06202623,
// 32'h06304103,
// 32'h06202823,
// 32'h06005103,
// 32'h06202a23,
// 32'h06105103,
// 32'h06202c23,
// 32'h06205103,
// 32'h06202e23,
// 32'h06305103,
// 32'h08202023,
// 32'haa0bc0b7,
// 32'h0dd08093,
// 32'h06102023,
// 32'h07700113,
// 32'h062001a3,
// 32'h06002183,
// 32'h06302223,
// 32'h01100113,
// 32'h06200123,
// 32'h06002183,
// 32'h06302423,
// 32'h02200113,
// 32'h062000a3,
// 32'h06002183,
// 32'h06302623,
// 32'h03300113,
// 32'h06200023,
// 32'h06002183,
// 32'h06302823,
// 32'haa0bc0b7,
// 32'h0dd08093,
// 32'h06102023,
// 32'h0aa00113,
// 32'h00811113,
// 32'h0bb10113,
// 32'h062011a3,
// 32'h06002183,
// 32'h06302a23,
// 32'h0cc00113,
// 32'h00811113,
// 32'h0dd10113,
// 32'h06201123,
// 32'h06002183,
// 32'h06302c23,
// 32'h03300113,
// 32'h00811113,
// 32'h04410113,
// 32'h062010a3,
// 32'h06002183,
// 32'h06302e23,
// 32'h05500113,
// 32'h00811113,
// 32'h06610113,
// 32'h06201023,
// 32'h06002183,
// 32'h08302023,
// 32'h01e00113,
// 32'h02202423
//};